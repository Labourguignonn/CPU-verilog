module mult(
    input wire [31:0] A_in,
  	input wire [31:0] B_in, 
  	output reg [31:0] Hi,
  	output reg [31:0] Lo
    
);